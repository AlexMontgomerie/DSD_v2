module design_test_top;



endmodule