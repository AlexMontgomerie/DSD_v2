module ahfp_buf(in,
				out
				);
				
endmodule